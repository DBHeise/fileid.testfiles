version https://git-lfs.github.com/spec/v1
oid sha256:ac9734916562bd83aaa636f1746e49bd90ed15f9fd37f263acee7df4f3311a5c
size 16785408
